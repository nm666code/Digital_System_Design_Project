library verilog;
use verilog.vl_types.all;
entity motion_vlg_vec_tst is
end motion_vlg_vec_tst;
